bind game_fsm fsm_btn_interface_properties #(.ASSUME_MODE(1)) fsm_btn_interface_properties_i(.*);
